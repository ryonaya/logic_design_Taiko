module slide_pixel_decode(
    input  [2-1:0]  pre_slide_pixel,
    output [12-1:0] slide_pixel
);

parameter [12-1:0] list [0:3] = {
    12'h444,
    12'h666,
    12'h777,
    12'hBBB 
};
assign slide_pixel = list[pre_slide_pixel];

endmodule


module background_pixel_decode(
    input  [7-1:0]  pre_background_pixel,
    output [12-1:0] background_pixel
);

parameter [12-1:0] list [0:124] = {
    12'hFC8,
    12'hFE8,
    12'hEC8,
    12'hFE9,
    12'hFD8,
    12'h777,
    12'h000,
    12'h100,
    12'h332,
    12'hA87,
    12'hEB8,
    12'h925,
    12'hC26,
    12'h411,
    12'h211,
    12'h783,
    12'h711,
    12'hE27,
    12'h754,
    12'hC97,
    12'hFD7,
    12'h544,
    12'h666,
    12'hFEA,
    12'hFE6,
    12'hECA,
    12'hF9A,
    12'hCCB,
    12'hFEC,
    12'hFFF,
    12'hFCD,
    12'hFED,
    12'hFB7,
    12'hFDB,
    12'hF98,
    12'hC69,
    12'hDDD,
    12'hFC6,
    12'hCB9,
    12'hDB5,
    12'hBA4,
    12'hFD5,
    12'hFA6,
    12'hFCA,
    12'hFC5,
    12'hAAA,
    12'h998,
    12'hE7D,
    12'hE95,
    12'h642,
    12'h223,
    12'hFE4,
    12'h562,
    12'hFFD,
    12'hEB3,
    12'hDD3,
    12'hFB4,
    12'h333,
    12'hA74,
    12'hFC3,
    12'hDA2,
    12'hFD3,
    12'hFFC,
    12'hFFB,
    12'hCC3,
    12'h531,
    12'hD83,
    12'h962,
    12'hF84,
    12'hE92,
    12'hBEB,
    12'hFA3,
    12'hBC7,
    12'hDE8,
    12'hFB3,
    12'hDE5,
    12'hDEA,
    12'hEEE,
    12'hAB2,
    12'hB82,
    12'hFB2,
    12'hEFC,
    12'h852,
    12'hF94,
    12'hADD,
    12'hBEE,
    12'h8CD,
    12'h9EA,
    12'h5BD,
    12'h6BB,
    12'hFC0,
    12'h8ED,
    12'hF91,
    12'h7DA,
    12'hF61,
    12'hF82,
    12'hF72,
    12'hF63,
    12'h8A3,
    12'hD53,
    12'hA42,
    12'h9A2,
    12'h366,
    12'h478,
    12'h921,
    12'hDE1,
    12'hCD3,
    12'hBD3,
    12'h69A,
    12'hF93,
    12'h727,
    12'hB8F,
    12'h2D8,
    12'h3C3,
    12'h8C2,
    12'h97B,
    12'h3AB,
    12'hAD2,
    12'h425,
    12'hF52,
    12'hF74,
    12'hF42,
    12'hD10,
    12'hE21,
    12'hC20 
};
assign background_pixel = list[pre_background_pixel];

endmodule